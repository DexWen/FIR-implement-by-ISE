`timescale 1ms / 1us
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:53:39 03/30/2016 
// Design Name: 
// Module Name:    fix_mult 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fix_mult ( clk,rst_n,in_a,in_b,y_out ); //16??????????,??32??????

  input clk,rst_n;
  input [15:0]   in_a,in_b; //??16??????
  output[31:0]   y_out;     //??32??????

  reg[31:0]   y_out;         //????,?????????
  reg[15:0]   x1,x2,x3,x4;   //x1,x2????????;x3?x4???????????
  reg         x5;            //???????????
  reg[29:0]   x6;            //30????,??15?????????
  reg[31:0]   x7;            //???????????
 
 always@ (negedge clk )
	 begin
		if(!rst_n )              //????,?????
			begin
			x1<=16'b0;
			x2<=16'b0;
			x3<=16'b0;
			x4<=16'b0;
			x5<=1'b0;
			x6<=30'b0;
			x7<=32'b0;
			y_out<=32'b0;
			end
		else
			 begin
			 x1<=in_a;             //???????
			 x2<=in_b;
			 x3<=(x1[15]==0)?x1:{x1[15],~x1[14:0]+1'b1};     //????????1,?????????,?????????1,????????,??????????
			 x4<=(x2[15]==0)?x2:{x2[15],~x2[14:0]+1'b1};     //??
			 x5<=x3[15]^x4[15];                              //??????????,?????????
			 x6<=x3[14:0]*x4[14:0];                          //??15???????
			 x7<={x5,x6,1'b0};                               //????????,?1????,30???????1????0??,??32???
			 y_out<=(x7[31]==0)?x7:{x7[31],~x7[30:0]+1'b1};  //??????????,?????????????
			 end
	 end
endmodule
